/**********************************************
 * Jesus Luciano
 * 4/2/20
 *
 * TOP.v
 *
 * Top Level Module for Intel 8008
 *
 *
 *
 *
 **********************************************/
module TOP();






endmodule